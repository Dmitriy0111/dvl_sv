/*
*  File            :   dvv_vm_pkg.sv
*  Autor           :   Vlasov D.V.
*  Data            :   2019.12.25
*  Language        :   SystemVerilog
*  Description     :   This is dvv packet
*  Copyright(c)    :   2019 Vlasov D.V.
*/

package dvv_vm_pkg;
    
    `include "dvv_classes/dvv_cc.sv"

    `include "dvv_classes/dvv_bc.sv"

    `include "dvv_classes/dvv_res.sv"
    `include "dvv_classes/dvv_res_db.sv"
    
    `include "dvv_classes/dvv_sock.sv"

endpackage : dvv_vm_pkg
